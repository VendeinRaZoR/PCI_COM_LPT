library verilog;
use verilog.vl_types.all;
entity PCI_target_controller is
    generic(
        CS_RESET        : integer := 0;
        CS_IDLE         : integer := 1;
        CS_READ         : integer := 2;
        CS_VIDPID_WRITE_DEVICE0: integer := 18;
        CS_STATUSCOMMAND_WRITE_DEVICE0: integer := 19;
        CS_CLASSCODE_WRITE_DEVICE0: integer := 20;
        CS_BIST_HEADER_LAT_CACH_WRITE_DEVICE0: integer := 21;
        CS_BAR0_WRITE_DEVICE0: integer := 22;
        CS_BAR1_WRITE_DEVICE0: integer := 23;
        CS_BAR2_WRITE_DEVICE0: integer := 24;
        CS_BAR3_WRITE_DEVICE0: integer := 25;
        CS_BAR4_WRITE_DEVICE0: integer := 26;
        CS_BAR5_WRITE_DEVICE0: integer := 27;
        CS_CARDBUS_WRITE_DEVICE0: integer := 28;
        CS_SUBSYSTEM_VENDOR_WRITE_DEVICE0: integer := 29;
        CS_EXPANSION_ROM_BAR_WRITE_DEVICE0: integer := 30;
        CS_CAP_POINTER_WRITE_DEVICE0: integer := 31;
        CS_LAT_INTERRUPT_WRITE_DEVICE0: integer := 32;
        CS_VIDPID_WRITE_DEVICE1: integer := 50;
        CS_STATUSCOMMAND_WRITE_DEVICE1: integer := 51;
        CS_CLASSCODE_WRITE_DEVICE1: integer := 52;
        CS_BIST_HEADER_LAT_CACH_WRITE_DEVICE1: integer := 53;
        CS_BAR0_WRITE_DEVICE1: integer := 54;
        CS_BAR1_WRITE_DEVICE1: integer := 55;
        CS_BAR2_WRITE_DEVICE1: integer := 56;
        CS_BAR3_WRITE_DEVICE1: integer := 57;
        CS_BAR4_WRITE_DEVICE1: integer := 58;
        CS_BAR5_WRITE_DEVICE1: integer := 59;
        CS_CARDBUS_WRITE_DEVICE1: integer := 60;
        CS_SUBSYSTEM_VENDOR_WRITE_DEVICE1: integer := 61;
        CS_EXPANSION_ROM_BAR_WRITE_DEVICE1: integer := 62;
        CS_CAP_POINTER_WRITE_DEVICE1: integer := 63;
        CS_LAT_INTERRUPT_WRITE_DEVICE1: integer := 64;
        CS_NULL         : integer := 125;
        CS_RESERVED     : integer := 126;
        INT_PIN_DEVICE0 : integer := 512;
        INT_PIN_DEVICE1 : integer := 256;
        INT_PIN_DEVICE2 : integer := 768;
        INT_PIN_DEVICE3 : integer := 1024;
        STATUS_MASK_DEVICE0: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        STATUS_MASK_DEVICE1: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        STATUS_MASK_DEVICE2: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        STATUS_MASK_DEVICE3: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        COMMAND_MASK_DEVICE0: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        COMMAND_MASK_DEVICE1: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        COMMAND_MASK_DEVICE2: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        COMMAND_MASK_DEVICE3: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        TRDY_DELAY      : integer := 0;
        MULTIFUNCTIONAL_DEVICE0: integer := 8388608;
        MULTIFUNCTIONAL_DEVICE1: integer := 8388608;
        MULTIFUNCTIONAL_DEVICE2: integer := 8388608;
        MULTIFUNCTIONAL_DEVICE3: integer := 8388608;
        VIDPID_DEVICE0  : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1);
        CLASSCODE_DEVICE0: integer := 201523280;
        VIDPID_DEVICE1  : integer := 1347633992;
        CLASSCODE_DEVICE1: integer := 117441039;
        VIDPID_DEVICE2  : integer := 0;
        CLASSCODE_DEVICE2: integer := 0;
        VIDPID_DEVICE3  : integer := 0;
        CLASSCODE_DEVICE3: integer := 0
    );
    port(
        clk             : in     vl_logic;
        addr_data       : inout  vl_logic_vector(31 downto 0);
        cbe             : in     vl_logic_vector(3 downto 0);
        idsel           : in     vl_logic;
        frame           : in     vl_logic;
        irdy            : in     vl_logic;
        devsel          : inout  vl_logic;
        trdy            : inout  vl_logic;
        reset           : in     vl_logic;
        par             : out    vl_logic;
        in_addr_offset_w_io: out    vl_logic_vector(7 downto 0);
        out_add_data_cs : out    vl_logic_vector(31 downto 0);
        in_command      : out    vl_logic_vector(3 downto 0);
        addr_data_buf_in_byte: out    vl_logic_vector(7 downto 0);
        addr_data_buf_in_word: out    vl_logic_vector(16 downto 0);
        addr_data_buf_in_dword: out    vl_logic_vector(32 downto 0);
        BAR0_DEVICE0_configured: out    vl_logic;
        BAR1_DEVICE0_configured: out    vl_logic;
        BAR2_DEVICE0_configured: out    vl_logic;
        BAR3_DEVICE0_configured: out    vl_logic;
        BAR4_DEVICE0_configured: out    vl_logic;
        BAR5_DEVICE0_configured: out    vl_logic;
        BAR0_DEVICE1_configured: out    vl_logic;
        BAR1_DEVICE1_configured: out    vl_logic;
        BAR2_DEVICE1_configured: out    vl_logic;
        BAR3_DEVICE1_configured: out    vl_logic;
        BAR4_DEVICE1_configured: out    vl_logic;
        BAR5_DEVICE1_configured: out    vl_logic;
        BAR0_DEVICE2_configured: out    vl_logic;
        BAR1_DEVICE2_configured: out    vl_logic;
        BAR2_DEVICE2_configured: out    vl_logic;
        BAR3_DEVICE2_configured: out    vl_logic;
        BAR4_DEVICE2_configured: out    vl_logic;
        BAR5_DEVICE2_configured: out    vl_logic;
        BAR0_DEVICE3_configured: out    vl_logic;
        BAR1_DEVICE3_configured: out    vl_logic;
        BAR2_DEVICE3_configured: out    vl_logic;
        BAR3_DEVICE3_configured: out    vl_logic;
        BAR4_DEVICE3_configured: out    vl_logic;
        BAR5_DEVICE3_configured: out    vl_logic;
        control         : out    vl_logic;
        is_config_space : out    vl_logic;
        is_BAR0_DEVICE0_address: out    vl_logic;
        is_BAR1_DEVICE0_address: out    vl_logic;
        is_BAR2_DEVICE0_address: out    vl_logic;
        is_BAR3_DEVICE0_address: out    vl_logic;
        is_BAR4_DEVICE0_address: out    vl_logic;
        is_BAR5_DEVICE0_address: out    vl_logic;
        is_BAR0_DEVICE1_address: out    vl_logic;
        is_BAR1_DEVICE1_address: out    vl_logic;
        is_BAR2_DEVICE1_address: out    vl_logic;
        is_BAR3_DEVICE1_address: out    vl_logic;
        is_BAR4_DEVICE1_address: out    vl_logic;
        is_BAR5_DEVICE1_address: out    vl_logic;
        is_BAR0_DEVICE2_address: out    vl_logic;
        is_BAR1_DEVICE2_address: out    vl_logic;
        is_BAR2_DEVICE2_address: out    vl_logic;
        is_BAR3_DEVICE2_address: out    vl_logic;
        is_BAR4_DEVICE2_address: out    vl_logic;
        is_BAR5_DEVICE2_address: out    vl_logic;
        is_BAR0_DEVICE3_address: out    vl_logic;
        is_BAR1_DEVICE3_address: out    vl_logic;
        is_BAR2_DEVICE3_address: out    vl_logic;
        is_BAR3_DEVICE3_address: out    vl_logic;
        is_BAR4_DEVICE3_address: out    vl_logic;
        is_BAR5_DEVICE3_address: out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CS_RESET : constant is 1;
    attribute mti_svvh_generic_type of CS_IDLE : constant is 1;
    attribute mti_svvh_generic_type of CS_READ : constant is 1;
    attribute mti_svvh_generic_type of CS_VIDPID_WRITE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CS_STATUSCOMMAND_WRITE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CS_CLASSCODE_WRITE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CS_BIST_HEADER_LAT_CACH_WRITE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CS_BAR0_WRITE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CS_BAR1_WRITE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CS_BAR2_WRITE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CS_BAR3_WRITE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CS_BAR4_WRITE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CS_BAR5_WRITE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CS_CARDBUS_WRITE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CS_SUBSYSTEM_VENDOR_WRITE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CS_EXPANSION_ROM_BAR_WRITE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CS_CAP_POINTER_WRITE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CS_LAT_INTERRUPT_WRITE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CS_VIDPID_WRITE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CS_STATUSCOMMAND_WRITE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CS_CLASSCODE_WRITE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CS_BIST_HEADER_LAT_CACH_WRITE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CS_BAR0_WRITE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CS_BAR1_WRITE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CS_BAR2_WRITE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CS_BAR3_WRITE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CS_BAR4_WRITE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CS_BAR5_WRITE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CS_CARDBUS_WRITE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CS_SUBSYSTEM_VENDOR_WRITE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CS_EXPANSION_ROM_BAR_WRITE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CS_CAP_POINTER_WRITE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CS_LAT_INTERRUPT_WRITE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CS_NULL : constant is 1;
    attribute mti_svvh_generic_type of CS_RESERVED : constant is 1;
    attribute mti_svvh_generic_type of INT_PIN_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of INT_PIN_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of INT_PIN_DEVICE2 : constant is 1;
    attribute mti_svvh_generic_type of INT_PIN_DEVICE3 : constant is 1;
    attribute mti_svvh_generic_type of STATUS_MASK_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of STATUS_MASK_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of STATUS_MASK_DEVICE2 : constant is 1;
    attribute mti_svvh_generic_type of STATUS_MASK_DEVICE3 : constant is 1;
    attribute mti_svvh_generic_type of COMMAND_MASK_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of COMMAND_MASK_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of COMMAND_MASK_DEVICE2 : constant is 1;
    attribute mti_svvh_generic_type of COMMAND_MASK_DEVICE3 : constant is 1;
    attribute mti_svvh_generic_type of TRDY_DELAY : constant is 1;
    attribute mti_svvh_generic_type of MULTIFUNCTIONAL_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of MULTIFUNCTIONAL_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of MULTIFUNCTIONAL_DEVICE2 : constant is 1;
    attribute mti_svvh_generic_type of MULTIFUNCTIONAL_DEVICE3 : constant is 1;
    attribute mti_svvh_generic_type of VIDPID_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of CLASSCODE_DEVICE0 : constant is 1;
    attribute mti_svvh_generic_type of VIDPID_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of CLASSCODE_DEVICE1 : constant is 1;
    attribute mti_svvh_generic_type of VIDPID_DEVICE2 : constant is 1;
    attribute mti_svvh_generic_type of CLASSCODE_DEVICE2 : constant is 1;
    attribute mti_svvh_generic_type of VIDPID_DEVICE3 : constant is 1;
    attribute mti_svvh_generic_type of CLASSCODE_DEVICE3 : constant is 1;
end PCI_target_controller;
