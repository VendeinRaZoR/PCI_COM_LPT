library verilog;
use verilog.vl_types.all;
entity COM_controller_16C550 is
    generic(
        TRDY_DELAY      : integer := 0;
        COMF_RESET      : integer := 0;
        COMF_IDLE       : integer := 1;
        COMF_READ       : integer := 2;
        COMF_RX_READ    : integer := 3;
        COMF_TX_WRITE   : integer := 4;
        COMF_IER_WRITE  : integer := 5;
        COMF_IIR_WRITE  : integer := 6;
        COMF_FCR_WRITE  : integer := 7;
        COMF_LCR_WRITE  : integer := 8;
        COMF_MCR_WRITE  : integer := 9;
        COMF_LSR_WRITE  : integer := 10;
        COMF_MSR_WRITE  : integer := 11;
        COMF_SCR_WRITE  : integer := 12;
        COMF_DLL_WRITE  : integer := 13;
        COMF_DLM_WRITE  : integer := 14;
        COMF_DLL_READ   : integer := 15;
        COMF_DLM_READ   : integer := 16;
        COMF_IIR_READ   : integer := 17;
        COMF_MCR_READ   : integer := 18;
        COMF_LCR_READ   : integer := 19;
        COMF_LSR_READ   : integer := 20;
        COMF_MSR_READ   : integer := 21;
        COMF_IER_READ   : integer := 22;
        COMF_TX_INT_FLAG_RESET: integer := 23;
        COMF_FIFO_WRITE : integer := 24;
        COMF_IER_CHECK  : integer := 25;
        COMF_TSR_ENABLE : integer := 26;
        COMF_RX_END     : integer := 27;
        COMF_RX_INT_FLAG_RESET: integer := 28;
        COMF_MODEM_INT_FLAG_RESET: integer := 29;
        COMF_LINE_INT_FLAG_RESET: integer := 30;
        COMF_TX_END     : integer := 31
    );
    port(
        clk             : in     vl_logic;
        irdy            : in     vl_logic;
        reset           : in     vl_logic;
        baudclk_221184kHz: in     vl_logic;
        RX1             : in     vl_logic;
        CTS             : in     vl_logic;
        DSR             : in     vl_logic;
        RI              : in     vl_logic;
        DCD             : in     vl_logic;
        in_addr_bar_offset_w_io: in     vl_logic_vector(7 downto 0);
        is_COM_configured: in     vl_logic;
        is_COM_iospace  : in     vl_logic;
        addr_data_buf_in_byte: in     vl_logic_vector(7 downto 0);
        in_command      : in     vl_logic_vector(3 downto 0);
        devsel          : out    vl_logic;
        trdy            : out    vl_logic;
        par             : out    vl_logic;
        interrupt_pin   : out    vl_logic;
        TX1             : out    vl_logic;
        RTS             : out    vl_logic;
        DTR             : out    vl_logic;
        control         : out    vl_logic;
        out_add_data_io : out    vl_logic_vector(31 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of TRDY_DELAY : constant is 1;
    attribute mti_svvh_generic_type of COMF_RESET : constant is 1;
    attribute mti_svvh_generic_type of COMF_IDLE : constant is 1;
    attribute mti_svvh_generic_type of COMF_READ : constant is 1;
    attribute mti_svvh_generic_type of COMF_RX_READ : constant is 1;
    attribute mti_svvh_generic_type of COMF_TX_WRITE : constant is 1;
    attribute mti_svvh_generic_type of COMF_IER_WRITE : constant is 1;
    attribute mti_svvh_generic_type of COMF_IIR_WRITE : constant is 1;
    attribute mti_svvh_generic_type of COMF_FCR_WRITE : constant is 1;
    attribute mti_svvh_generic_type of COMF_LCR_WRITE : constant is 1;
    attribute mti_svvh_generic_type of COMF_MCR_WRITE : constant is 1;
    attribute mti_svvh_generic_type of COMF_LSR_WRITE : constant is 1;
    attribute mti_svvh_generic_type of COMF_MSR_WRITE : constant is 1;
    attribute mti_svvh_generic_type of COMF_SCR_WRITE : constant is 1;
    attribute mti_svvh_generic_type of COMF_DLL_WRITE : constant is 1;
    attribute mti_svvh_generic_type of COMF_DLM_WRITE : constant is 1;
    attribute mti_svvh_generic_type of COMF_DLL_READ : constant is 1;
    attribute mti_svvh_generic_type of COMF_DLM_READ : constant is 1;
    attribute mti_svvh_generic_type of COMF_IIR_READ : constant is 1;
    attribute mti_svvh_generic_type of COMF_MCR_READ : constant is 1;
    attribute mti_svvh_generic_type of COMF_LCR_READ : constant is 1;
    attribute mti_svvh_generic_type of COMF_LSR_READ : constant is 1;
    attribute mti_svvh_generic_type of COMF_MSR_READ : constant is 1;
    attribute mti_svvh_generic_type of COMF_IER_READ : constant is 1;
    attribute mti_svvh_generic_type of COMF_TX_INT_FLAG_RESET : constant is 1;
    attribute mti_svvh_generic_type of COMF_FIFO_WRITE : constant is 1;
    attribute mti_svvh_generic_type of COMF_IER_CHECK : constant is 1;
    attribute mti_svvh_generic_type of COMF_TSR_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of COMF_RX_END : constant is 1;
    attribute mti_svvh_generic_type of COMF_RX_INT_FLAG_RESET : constant is 1;
    attribute mti_svvh_generic_type of COMF_MODEM_INT_FLAG_RESET : constant is 1;
    attribute mti_svvh_generic_type of COMF_LINE_INT_FLAG_RESET : constant is 1;
    attribute mti_svvh_generic_type of COMF_TX_END : constant is 1;
end COM_controller_16C550;
