library verilog;
use verilog.vl_types.all;
entity pci_com_lpt_usb_eth_vlg_tst is
end pci_com_lpt_usb_eth_vlg_tst;
